`include "mips_defines.v"

module cache (
    input clk,
    input memclk,
    input [31:0] addr, // byte address
    input we,
    input re,
    input rst,
    input [31:0] din,

    output wire [31:0] dout,
    output wire complete
);

    // when implementing your cache FSM logic
    // you will write and read from these structures
    // containing the valid bits, tag, and data, for each cache
    // block, indexed from 0 to 63
    // you may modify these structures to implement more complicated caches,
    // but their total size must not increase

    // this will support 64 blocks of 4 words each, for a total of 1KB of
    // cache data storage
    reg valid_bits [63:0];
    reg [21:0] tag_bits [63:0];
    reg [127:0] data_blocks [63:0];

    // outputs from DRAM
    wire [127:0] dram_out;
    wire dram_complete;

    // USE THIS SYNCHRONOUS BLOCK TO ASSIGN THE INPUTS TO DRAM
    
    // inputs to dram should be regs when assigned in a state machine
    reg dram_we, dram_re;
    wire [`MEM_DEPTH-3:0] dram_addr = {addr[`MEM_DEPTH-1:4], 2'b0};  
		// *** ??? this would get to the beginning of that block (minus the block offset) + 2b'0 --> i.e. beginning of the block instead of word in the block's address?
    reg [127:0] dram_in;
    reg [31:0] cache_dout;
    reg cache_complete;
    wire [5:0] index = addr[9:4];
    reg [127:0] block;
    wire [1:0] block_start = addr[3:2];

	integer i;
	initial begin
		for (i = 0; i <= 63; i = i+1) begin
			valid_bits [i] = 1'b0;
			tag_bits [i] = 22'b0;
			data_blocks [i] = 128'b0;
		end
	end

    /* Need to account for:
     * re 
     *   - compulsory miss
     *   - conflict miss
     *      dram -> cache
     *      cache -> dout
     *   - hit
     *      cache -> dout
     * we
     *   - miss
     *      din -> dram
     *   - hit
     *      din -> cache
     *      din -> dram
     */

    //determine whether or not input is in cache
    // index = addr[8:4]
    // is valid_bits[index] == 1?
    // is tag_bits == addr[31:8]
    wire cache_hit = (valid_bits[index] == 1'b1) && (tag_bits[index] == addr[31:10]); 

    always @(posedge clk or negedge rst) begin
	if (~rst) begin
	    dram_in <= 128'b0;
	    cache_dout <= 32'b0;
	    cache_complete <= 1'b1;
	    block <= 128'b0;
	end
        // if (re)  //reading
        if ( re == 1'b1 ) begin
            //dram_we = 1b'0;
            dram_we <= 1'b0;
            //not in cache // (miss)
            if ( cache_hit == 1'b0 ) begin
                dram_re <= 1'b1;
                //set cache
                    valid_bits[index] <= 1;
                    tag_bits[index] <= addr[31:10];
                    data_blocks[index] <= dram_out;
                cache_dout <= dram_out;
                cache_complete <= dram_complete;
            end
				
            //in cache // (hit)
            if ( cache_hit == 1'b1 ) begin
                dram_re = 1'b0;
                //calc cache_dout
                    block = data_blocks[index];
                    case (block_start)
                        2'b00: cache_dout = block[31:0];
                        2'b01: cache_dout = block[63:32];
                        2'b10: cache_dout = block[95:64];
                        2'b11: cache_dout = block[127:96];
                    endcase
                cache_complete = ~ (re | we);  //***???
            end
				
        end
        // if (we)
        if ( we == 1'b1 ) begin    
            dram_re = 1'b0;
			dram_we = 1'b1;
            //not in cache  // (miss) --> 
			if ( cache_hit == 1'b0 ) begin
                //dram_in[block_start + 31: block_start] = din;
                case (block_start)
                    2'b00: dram_in[31:0] = din;
                    2'b01: dram_in[63:32] = din;
                    2'b10: dram_in[95:64] = din;
                    2'b11: dram_in[127:96] = din;
                endcase
                cache_complete = dram_complete;
			end
				
            //in cache  // (hit)
			if ( cache_hit == 1'b1 ) begin
               // dram_in[block_start + 31: block_start] = din;
                //set cache
                    //index = addr[8:4]
					block = data_blocks[index];
                    //block [block_start + 31: block_start] = din;
                case (block_start)
                    2'b00: begin
                        data_blocks[index][31:0] = din;
                        dram_in[31:0] = din;
                    end
                    2'b01: begin
                        data_blocks[index][63:32] = din;
                        dram_in[63:32] = din;
                    end
                    2'b10: begin
                        data_blocks[index][95:64] = din;
                        dram_in[95:64] = din;
                    end
                    2'b11: begin
                        data_blocks[index][127:96] = din;
                        dram_in[127:96] = din;
                    end
                endcase
                cache_complete = dram_complete;
			end
                
        end

    end
    
    

    // COMMENT OUT THIS CONTINUOUS CODE WHEN IMPLEMENTING YOUR CACHE
    // The code below implements the cache module in the trivial case when
    // we don't use a cache and we use only the first word in each memory
    // block, (which are four words each).
    /*

    // just pass we and re straignt to the DRAM
    wire dram_we = we;
    wire dram_re = re;

    // address a whole block per word (2^4 bytes)
    // change this in your implementation
    wire [`MEM_DEPTH-3:0] dram_addr = addr[`MEM_DEPTH-1:2];

    // only use the first word in the cache line
    // change this in your implementation
    wire [127:0] dram_in = {96'd0, din};
    wire [31:0] cache_dout = dram_out[31:0];

    // the cache is done when DRAM is done
    wire cache_complete = dram_complete;

    */

    dataram dram (.clk(clk),
                  .memclk(memclk),
                  .rst(rst),
                  .we(dram_we),
                  .re(dram_re),
                  .addr(dram_addr),
                  .din(dram_in),
                  .dout(dram_out),
                  .complete(dram_complete));
    
    assign dout = cache_dout;
    assign complete = cache_complete;

endmodule
