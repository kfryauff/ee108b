// Custom IROM with self-playing Pong

`include "mips_defines.v"

`define ADDR_WIDTH 9
`define INSTR_WIDTH 32
`define NUM_INSTR 512

module irom(addr, dout);
  input [`ADDR_WIDTH-1:0] addr;
  output wire [`INSTR_WIDTH-1:0] dout;

  wire [`INSTR_WIDTH-1:0] memory [`NUM_INSTR-1:0];

  assign dout = memory[addr];

assign memory[0] = {`ORI, `ZERO, `T0, 16'hffff};
assign memory[1] = {`ANDI, `ZERO, `T1, 16'd0};

assign memory[2]={`SW, `T1, `T0, 16'd2312};

assign memory[4]={`SW, `T1, `T0, 16'd884};

assign memory[6]={`SW, `T1, `T0, 16'd3688};

assign memory[8]={`SW, `T1, `T0, 16'd960};

assign memory[10]={`SW, `T1, `T0, 16'd3416};

assign memory[12]={`SW, `T1, `T0, 16'd720};

assign memory[14]={`SW, `T1, `T0, 16'd2252};

assign memory[16]={`SW, `T1, `T0, 16'd2192};

assign memory[18]={`SW, `T1, `T0, 16'd1656};

assign memory[20]={`SW, `T1, `T0, 16'd2808};

assign memory[22]={`SW, `T1, `T0, 16'd3600};

assign memory[24]={`SW, `T1, `T0, 16'd1108};

assign memory[26]={`SW, `T1, `T0, 16'd3204};

assign memory[28]={`SW, `T1, `T0, 16'd2676};

assign memory[30]={`SW, `T1, `T0, 16'd3252};

assign memory[32]={`SW, `T1, `T0, 16'd3920};

assign memory[34]={`SW, `T1, `T0, 16'd3384};

assign memory[36]={`SW, `T1, `T0, 16'd1108};

assign memory[38]={`SW, `T1, `T0, 16'd3432};

assign memory[40]={`SW, `T1, `T0, 16'd1940};

assign memory[42]={`SW, `T1, `T0, 16'd728};

assign memory[44]={`SW, `T1, `T0, 16'd684};

assign memory[46]={`SW, `T1, `T0, 16'd3952};

assign memory[48]={`SW, `T1, `T0, 16'd2760};

assign memory[50]={`SW, `T1, `T0, 16'd2308};

assign memory[52]={`SW, `T1, `T0, 16'd3432};

assign memory[54]={`SW, `T1, `T0, 16'd3560};

assign memory[56]={`SW, `T1, `T0, 16'd1232};

assign memory[58]={`SW, `T1, `T0, 16'd2288};

assign memory[60]={`SW, `T1, `T0, 16'd3336};

assign memory[62]={`SW, `T1, `T0, 16'd112};

assign memory[64]={`SW, `T1, `T0, 16'd2252};

assign memory[66]={`SW, `T1, `T0, 16'd3116};

assign memory[68]={`SW, `T1, `T0, 16'd12};

assign memory[70]={`SW, `T1, `T0, 16'd2052};

assign memory[72]={`SW, `T1, `T0, 16'd916};

assign memory[74]={`SW, `T1, `T0, 16'd2752};

assign memory[76]={`SW, `T1, `T0, 16'd2304};

assign memory[78]={`SW, `T1, `T0, 16'd3640};

assign memory[80]={`SW, `T1, `T0, 16'd3344};

assign memory[82]={`SW, `T1, `T0, 16'd816};

assign memory[84]={`SW, `T1, `T0, 16'd2692};

assign memory[86]={`SW, `T1, `T0, 16'd2364};

assign memory[88]={`SW, `T1, `T0, 16'd2136};

assign memory[90]={`SW, `T1, `T0, 16'd780};

assign memory[92]={`SW, `T1, `T0, 16'd344};

assign memory[94]={`SW, `T1, `T0, 16'd2744};

assign memory[96]={`SW, `T1, `T0, 16'd632};

assign memory[98]={`SW, `T1, `T0, 16'd2748};

assign memory[100]={`SW, `T1, `T0, 16'd3712};

assign memory[102]={`SW, `T1, `T0, 16'd12};

assign memory[104]={`SW, `T1, `T0, 16'd212};

assign memory[106]={`SW, `T1, `T0, 16'd2928};

assign memory[108]={`SW, `T1, `T0, 16'd808};

assign memory[110]={`SW, `T1, `T0, 16'd3420};

assign memory[112]={`SW, `T1, `T0, 16'd1000};

assign memory[114]={`SW, `T1, `T0, 16'd2028};

assign memory[116]={`SW, `T1, `T0, 16'd1180};

assign memory[118]={`SW, `T1, `T0, 16'd3060};

assign memory[120]={`SW, `T1, `T0, 16'd1528};

assign memory[122]={`SW, `T1, `T0, 16'd1164};

assign memory[124]={`SW, `T1, `T0, 16'd1960};

assign memory[126]={`SW, `T1, `T0, 16'd2380};

assign memory[128]={`SW, `T1, `T0, 16'd2528};

assign memory[130]={`SW, `T1, `T0, 16'd1704};

assign memory[132]={`SW, `T1, `T0, 16'd60};

assign memory[134]={`SW, `T1, `T0, 16'd304};

assign memory[136]={`SW, `T1, `T0, 16'd1244};

assign memory[138]={`SW, `T1, `T0, 16'd1144};

assign memory[140]={`SW, `T1, `T0, 16'd1352};

assign memory[142]={`SW, `T1, `T0, 16'd3244};

assign memory[144]={`SW, `T1, `T0, 16'd3660};

assign memory[146]={`SW, `T1, `T0, 16'd236};

assign memory[148]={`SW, `T1, `T0, 16'd3084};

assign memory[150]={`SW, `T1, `T0, 16'd376};

assign memory[152]={`SW, `T1, `T0, 16'd3120};

assign memory[154]={`SW, `T1, `T0, 16'd1792};

assign memory[156]={`SW, `T1, `T0, 16'd428};

assign memory[158]={`SW, `T1, `T0, 16'd3800};

assign memory[160]={`SW, `T1, `T0, 16'd3276};

assign memory[162]={`SW, `T1, `T0, 16'd160};

assign memory[164]={`SW, `T1, `T0, 16'd196};

assign memory[166]={`SW, `T1, `T0, 16'd436};

assign memory[168]={`SW, `T1, `T0, 16'd2452};

assign memory[170]={`SW, `T1, `T0, 16'd3328};

assign memory[172]={`SW, `T1, `T0, 16'd96};

assign memory[174]={`SW, `T1, `T0, 16'd3012};

assign memory[176]={`SW, `T1, `T0, 16'd2856};

assign memory[178]={`SW, `T1, `T0, 16'd3356};

assign memory[180]={`SW, `T1, `T0, 16'd572};

assign memory[182]={`SW, `T1, `T0, 16'd3688};

assign memory[184]={`SW, `T1, `T0, 16'd128};

assign memory[186]={`SW, `T1, `T0, 16'd3264};

assign memory[188]={`SW, `T1, `T0, 16'd3004};

assign memory[190]={`SW, `T1, `T0, 16'd3824};

assign memory[192]={`SW, `T1, `T0, 16'd3988};

assign memory[194]={`SW, `T1, `T0, 16'd2308};

assign memory[196]={`SW, `T1, `T0, 16'd2996};

assign memory[198]={`SW, `T1, `T0, 16'd1900};

assign memory[200]={`SW, `T1, `T0, 16'd1844};

assign memory[202]={`SW, `T1, `T0, 16'd2952};

assign memory[204]={`SW, `T1, `T0, 16'd572};

assign memory[206]={`SW, `T1, `T0, 16'd2588};

assign memory[208]={`SW, `T1, `T0, 16'd2908};

assign memory[210]={`SW, `T1, `T0, 16'd3116};

assign memory[212]={`SW, `T1, `T0, 16'd944};

assign memory[214]={`SW, `T1, `T0, 16'd3528};

assign memory[216]={`SW, `T1, `T0, 16'd208};

assign memory[218]={`SW, `T1, `T0, 16'd3704};

assign memory[220]={`SW, `T1, `T0, 16'd2920};

assign memory[222]={`SW, `T1, `T0, 16'd3700};

assign memory[224]={`SW, `T1, `T0, 16'd3192};

assign memory[226]={`SW, `T1, `T0, 16'd1788};

assign memory[228]={`SW, `T1, `T0, 16'd272};

assign memory[230]={`SW, `T1, `T0, 16'd3004};

assign memory[232]={`SW, `T1, `T0, 16'd3464};

assign memory[234]={`SW, `T1, `T0, 16'd3892};

assign memory[236]={`SW, `T1, `T0, 16'd1952};

assign memory[238]={`SW, `T1, `T0, 16'd1344};

assign memory[240]={`SW, `T1, `T0, 16'd1116};

assign memory[242]={`SW, `T1, `T0, 16'd4056};

assign memory[244]={`SW, `T1, `T0, 16'd540};

assign memory[246]={`SW, `T1, `T0, 16'd416};

assign memory[248]={`SW, `T1, `T0, 16'd564};

assign memory[250]={`SW, `T1, `T0, 16'd1596};

assign memory[252]={`SW, `T1, `T0, 16'd3640};

assign memory[254]={`SW, `T1, `T0, 16'd624};

assign memory[256]={`SW, `T1, `T0, 16'd3380};

assign memory[258]={`SW, `T1, `T0, 16'd2672};

assign memory[260]={`SW, `T1, `T0, 16'd820};

assign memory[262]={`SW, `T1, `T0, 16'd2496};

assign memory[264]={`SW, `T1, `T0, 16'd892};

assign memory[266]={`SW, `T1, `T0, 16'd584};

assign memory[268]={`SW, `T1, `T0, 16'd264};

assign memory[270]={`SW, `T1, `T0, 16'd156};

assign memory[272]={`SW, `T1, `T0, 16'd412};

assign memory[274]={`SW, `T1, `T0, 16'd2484};

assign memory[276]={`SW, `T1, `T0, 16'd3192};

assign memory[278]={`SW, `T1, `T0, 16'd64};

assign memory[280]={`SW, `T1, `T0, 16'd3888};

assign memory[282]={`SW, `T1, `T0, 16'd1944};

assign memory[284]={`SW, `T1, `T0, 16'd1540};

assign memory[286]={`SW, `T1, `T0, 16'd1188};

assign memory[288]={`SW, `T1, `T0, 16'd2712};

assign memory[290]={`SW, `T1, `T0, 16'd2204};

assign memory[292]={`SW, `T1, `T0, 16'd2136};

assign memory[294]={`SW, `T1, `T0, 16'd2808};

assign memory[296]={`SW, `T1, `T0, 16'd3340};

assign memory[298]={`SW, `T1, `T0, 16'd1100};

assign memory[300]={`SW, `T1, `T0, 16'd2272};

assign memory[302]={`SW, `T1, `T0, 16'd3796};

assign memory[304]={`SW, `T1, `T0, 16'd1840};

assign memory[306]={`SW, `T1, `T0, 16'd268};

assign memory[308]={`SW, `T1, `T0, 16'd76};

assign memory[310]={`SW, `T1, `T0, 16'd476};

assign memory[312]={`SW, `T1, `T0, 16'd2476};

assign memory[314]={`SW, `T1, `T0, 16'd1272};

assign memory[316]={`SW, `T1, `T0, 16'd3748};

assign memory[318]={`SW, `T1, `T0, 16'd3264};

assign memory[320]={`SW, `T1, `T0, 16'd1564};

assign memory[322]={`SW, `T1, `T0, 16'd1440};

assign memory[324]={`SW, `T1, `T0, 16'd3152};

assign memory[326]={`SW, `T1, `T0, 16'd496};

assign memory[328]={`SW, `T1, `T0, 16'd3252};

assign memory[330]={`SW, `T1, `T0, 16'd3384};

assign memory[332]={`SW, `T1, `T0, 16'd256};

assign memory[334]={`SW, `T1, `T0, 16'd3556};

assign memory[336]={`SW, `T1, `T0, 16'd1824};

assign memory[338]={`SW, `T1, `T0, 16'd1412};

assign memory[340]={`SW, `T1, `T0, 16'd3152};

assign memory[342]={`SW, `T1, `T0, 16'd948};

assign memory[344]={`SW, `T1, `T0, 16'd2204};

assign memory[346]={`SW, `T1, `T0, 16'd2708};

assign memory[348]={`SW, `T1, `T0, 16'd2512};

assign memory[350]={`SW, `T1, `T0, 16'd2316};

assign memory[352]={`SW, `T1, `T0, 16'd1156};

assign memory[354]={`SW, `T1, `T0, 16'd2604};

assign memory[356]={`SW, `T1, `T0, 16'd2504};

assign memory[358]={`SW, `T1, `T0, 16'd2072};

assign memory[360]={`SW, `T1, `T0, 16'd2412};

assign memory[362]={`SW, `T1, `T0, 16'd1648};

assign memory[364]={`SW, `T1, `T0, 16'd3704};

assign memory[366]={`SW, `T1, `T0, 16'd252};

assign memory[368]={`SW, `T1, `T0, 16'd2008};

assign memory[370]={`SW, `T1, `T0, 16'd340};

assign memory[372]={`SW, `T1, `T0, 16'd1596};

assign memory[374]={`SW, `T1, `T0, 16'd3988};

assign memory[376]={`SW, `T1, `T0, 16'd1028};

assign memory[378]={`SW, `T1, `T0, 16'd3860};

assign memory[380]={`SW, `T1, `T0, 16'd496};

assign memory[382]={`SW, `T1, `T0, 16'd2220};

assign memory[384]={`SW, `T1, `T0, 16'd3132};

assign memory[386]={`SW, `T1, `T0, 16'd3276};

assign memory[388]={`SW, `T1, `T0, 16'd3376};

assign memory[390]={`SW, `T1, `T0, 16'd768};

assign memory[392]={`SW, `T1, `T0, 16'd2084};

assign memory[394]={`SW, `T1, `T0, 16'd892};

assign memory[396]={`SW, `T1, `T0, 16'd2588};

assign memory[398]={`SW, `T1, `T0, 16'd3404};

assign memory[400]={`SW, `T1, `T0, 16'd1948};

assign memory[402]={`SW, `T1, `T0, 16'd3380};

assign memory[404]={`SW, `T1, `T0, 16'd124};

assign memory[406]={`SW, `T1, `T0, 16'd1444};

assign memory[408]={`SW, `T1, `T0, 16'd116};

assign memory[410]={`SW, `T1, `T0, 16'd1808};

assign memory[412]={`SW, `T1, `T0, 16'd560};

assign memory[414]={`SW, `T1, `T0, 16'd3472};

assign memory[416]={`SW, `T1, `T0, 16'd1720};

assign memory[418]={`SW, `T1, `T0, 16'd568};

assign memory[420]={`SW, `T1, `T0, 16'd388};

assign memory[422]={`SW, `T1, `T0, 16'd1472};

assign memory[424]={`SW, `T1, `T0, 16'd2548};

assign memory[426]={`SW, `T1, `T0, 16'd3492};

assign memory[428]={`SW, `T1, `T0, 16'd108};

assign memory[430]={`SW, `T1, `T0, 16'd800};

assign memory[432]={`SW, `T1, `T0, 16'd2328};

assign memory[434]={`SW, `T1, `T0, 16'd640};

assign memory[436]={`SW, `T1, `T0, 16'd1076};

assign memory[438]={`SW, `T1, `T0, 16'd464};

assign memory[440]={`SW, `T1, `T0, 16'd2412};

assign memory[442]={`SW, `T1, `T0, 16'd1752};

assign memory[444]={`SW, `T1, `T0, 16'd528};

assign memory[446]={`SW, `T1, `T0, 16'd2576};

assign memory[448]={`SW, `T1, `T0, 16'd2944};

assign memory[450]={`SW, `T1, `T0, 16'd3192};

assign memory[452]={`SW, `T1, `T0, 16'd3776};

assign memory[454]={`SW, `T1, `T0, 16'd3072};

assign memory[456]={`SW, `T1, `T0, 16'd4028};

assign memory[458]={`SW, `T1, `T0, 16'd2404};

assign memory[460]={`SW, `T1, `T0, 16'd3240};

assign memory[462]={`SW, `T1, `T0, 16'd244};

assign memory[464]={`SW, `T1, `T0, 16'd3784};

assign memory[466]={`SW, `T1, `T0, 16'd2016};

assign memory[468]={`SW, `T1, `T0, 16'd3512};

assign memory[470]={`SW, `T1, `T0, 16'd3052};

assign memory[472]={`SW, `T1, `T0, 16'd2160};

assign memory[474]={`SW, `T1, `T0, 16'd3568};

assign memory[476]={`SW, `T1, `T0, 16'd456};

assign memory[478]={`SW, `T1, `T0, 16'd892};

assign memory[480]={`SW, `T1, `T0, 16'd3764};

assign memory[482]={`SW, `T1, `T0, 16'd4076};

assign memory[484]={`SW, `T1, `T0, 16'd3552};

assign memory[486]={`SW, `T1, `T0, 16'd564};

assign memory[488]={`SW, `T1, `T0, 16'd3924};

assign memory[490]={`SW, `T1, `T0, 16'd1984};

assign memory[492]={`SW, `T1, `T0, 16'd2512};

assign memory[494]={`SW, `T1, `T0, 16'd2140};

assign memory[496]={`SW, `T1, `T0, 16'd160};

assign memory[498]={`SW, `T1, `T0, 16'd1384};

assign memory[500]={`SW, `T1, `T0, 16'd80};

assign memory[502]={`SW, `T1, `T0, 16'd1656};

assign memory[504]={`SW, `T1, `T0, 16'd1356};

assign memory[506]={`SW, `T1, `T0, 16'd2252};

assign memory[508]={`SW, `T1, `T0, 16'd3824};

assign memory[510]={`SW, `T1, `T0, 16'd3988};

 assign memory[3]={`LW, `T1, `T0, 16'd2312};

assign memory[5]={`LW, `T1, `T0, 16'd884};

assign memory[7]={`LW, `T1, `T0, 16'd3688};

assign memory[9]={`LW, `T1, `T0, 16'd960};

assign memory[11]={`LW, `T1, `T0, 16'd3416};

assign memory[13]={`LW, `T1, `T0, 16'd720};

assign memory[15]={`LW, `T1, `T0, 16'd2252};

assign memory[17]={`LW, `T1, `T0, 16'd2192};

assign memory[19]={`LW, `T1, `T0, 16'd1656};

assign memory[21]={`LW, `T1, `T0, 16'd2808};

assign memory[23]={`LW, `T1, `T0, 16'd3600};

assign memory[25]={`LW, `T1, `T0, 16'd1108};

assign memory[27]={`LW, `T1, `T0, 16'd3204};

assign memory[29]={`LW, `T1, `T0, 16'd2676};

assign memory[31]={`LW, `T1, `T0, 16'd3252};

assign memory[33]={`LW, `T1, `T0, 16'd3920};

assign memory[35]={`LW, `T1, `T0, 16'd3384};

assign memory[37]={`LW, `T1, `T0, 16'd1108};

assign memory[39]={`LW, `T1, `T0, 16'd3432};

assign memory[41]={`LW, `T1, `T0, 16'd1940};

assign memory[43]={`LW, `T1, `T0, 16'd728};

assign memory[45]={`LW, `T1, `T0, 16'd684};

assign memory[47]={`LW, `T1, `T0, 16'd3952};

assign memory[49]={`LW, `T1, `T0, 16'd2760};

assign memory[51]={`LW, `T1, `T0, 16'd2308};

assign memory[53]={`LW, `T1, `T0, 16'd3432};

assign memory[55]={`LW, `T1, `T0, 16'd3560};

assign memory[57]={`LW, `T1, `T0, 16'd1232};

assign memory[59]={`LW, `T1, `T0, 16'd2288};

assign memory[61]={`LW, `T1, `T0, 16'd3336};

assign memory[63]={`LW, `T1, `T0, 16'd112};

assign memory[65]={`LW, `T1, `T0, 16'd2252};

assign memory[67]={`LW, `T1, `T0, 16'd3116};

assign memory[69]={`LW, `T1, `T0, 16'd12};

assign memory[71]={`LW, `T1, `T0, 16'd2052};

assign memory[73]={`LW, `T1, `T0, 16'd916};

assign memory[75]={`LW, `T1, `T0, 16'd2752};

assign memory[77]={`LW, `T1, `T0, 16'd2304};

assign memory[79]={`LW, `T1, `T0, 16'd3640};

assign memory[81]={`LW, `T1, `T0, 16'd3344};

assign memory[83]={`LW, `T1, `T0, 16'd816};

assign memory[85]={`LW, `T1, `T0, 16'd2692};

assign memory[87]={`LW, `T1, `T0, 16'd2364};

assign memory[89]={`LW, `T1, `T0, 16'd2136};

assign memory[91]={`LW, `T1, `T0, 16'd780};

assign memory[93]={`LW, `T1, `T0, 16'd344};

assign memory[95]={`LW, `T1, `T0, 16'd2744};

assign memory[97]={`LW, `T1, `T0, 16'd632};

assign memory[99]={`LW, `T1, `T0, 16'd2748};

assign memory[101]={`LW, `T1, `T0, 16'd3712};

assign memory[103]={`LW, `T1, `T0, 16'd12};

assign memory[105]={`LW, `T1, `T0, 16'd212};

assign memory[107]={`LW, `T1, `T0, 16'd2928};

assign memory[109]={`LW, `T1, `T0, 16'd808};

assign memory[111]={`LW, `T1, `T0, 16'd3420};

assign memory[113]={`LW, `T1, `T0, 16'd1000};

assign memory[115]={`LW, `T1, `T0, 16'd2028};

assign memory[117]={`LW, `T1, `T0, 16'd1180};

assign memory[119]={`LW, `T1, `T0, 16'd3060};

assign memory[121]={`LW, `T1, `T0, 16'd1528};

assign memory[123]={`LW, `T1, `T0, 16'd1164};

assign memory[125]={`LW, `T1, `T0, 16'd1960};

assign memory[127]={`LW, `T1, `T0, 16'd2380};

assign memory[129]={`LW, `T1, `T0, 16'd2528};

assign memory[131]={`LW, `T1, `T0, 16'd1704};

assign memory[133]={`LW, `T1, `T0, 16'd60};

assign memory[135]={`LW, `T1, `T0, 16'd304};

assign memory[137]={`LW, `T1, `T0, 16'd1244};

assign memory[139]={`LW, `T1, `T0, 16'd1144};

assign memory[141]={`LW, `T1, `T0, 16'd1352};

assign memory[143]={`LW, `T1, `T0, 16'd3244};

assign memory[145]={`LW, `T1, `T0, 16'd3660};

assign memory[147]={`LW, `T1, `T0, 16'd236};

assign memory[149]={`LW, `T1, `T0, 16'd3084};

assign memory[151]={`LW, `T1, `T0, 16'd376};

assign memory[153]={`LW, `T1, `T0, 16'd3120};

assign memory[155]={`LW, `T1, `T0, 16'd1792};

assign memory[157]={`LW, `T1, `T0, 16'd428};

assign memory[159]={`LW, `T1, `T0, 16'd3800};

assign memory[161]={`LW, `T1, `T0, 16'd3276};

assign memory[163]={`LW, `T1, `T0, 16'd160};

assign memory[165]={`LW, `T1, `T0, 16'd196};

assign memory[167]={`LW, `T1, `T0, 16'd436};

assign memory[169]={`LW, `T1, `T0, 16'd2452};

assign memory[171]={`LW, `T1, `T0, 16'd3328};

assign memory[173]={`LW, `T1, `T0, 16'd96};

assign memory[175]={`LW, `T1, `T0, 16'd3012};

assign memory[177]={`LW, `T1, `T0, 16'd2856};

assign memory[179]={`LW, `T1, `T0, 16'd3356};

assign memory[181]={`LW, `T1, `T0, 16'd572};

assign memory[183]={`LW, `T1, `T0, 16'd3688};

assign memory[185]={`LW, `T1, `T0, 16'd128};

assign memory[187]={`LW, `T1, `T0, 16'd3264};

assign memory[189]={`LW, `T1, `T0, 16'd3004};

assign memory[191]={`LW, `T1, `T0, 16'd3824};

assign memory[193]={`LW, `T1, `T0, 16'd3988};

assign memory[195]={`LW, `T1, `T0, 16'd2308};

assign memory[197]={`LW, `T1, `T0, 16'd2996};

assign memory[199]={`LW, `T1, `T0, 16'd1900};

assign memory[201]={`LW, `T1, `T0, 16'd1844};

assign memory[203]={`LW, `T1, `T0, 16'd2952};

assign memory[205]={`LW, `T1, `T0, 16'd572};

assign memory[207]={`LW, `T1, `T0, 16'd2588};

assign memory[209]={`LW, `T1, `T0, 16'd2908};

assign memory[211]={`LW, `T1, `T0, 16'd3116};

assign memory[213]={`LW, `T1, `T0, 16'd944};

assign memory[215]={`LW, `T1, `T0, 16'd3528};

assign memory[217]={`LW, `T1, `T0, 16'd208};

assign memory[219]={`LW, `T1, `T0, 16'd3704};

assign memory[221]={`LW, `T1, `T0, 16'd2920};

assign memory[223]={`LW, `T1, `T0, 16'd3700};

assign memory[225]={`LW, `T1, `T0, 16'd3192};

assign memory[227]={`LW, `T1, `T0, 16'd1788};

assign memory[229]={`LW, `T1, `T0, 16'd272};

assign memory[231]={`LW, `T1, `T0, 16'd3004};

assign memory[233]={`LW, `T1, `T0, 16'd3464};

assign memory[235]={`LW, `T1, `T0, 16'd3892};

assign memory[237]={`LW, `T1, `T0, 16'd1952};

assign memory[239]={`LW, `T1, `T0, 16'd1344};

assign memory[241]={`LW, `T1, `T0, 16'd1116};

assign memory[243]={`LW, `T1, `T0, 16'd4056};

assign memory[245]={`LW, `T1, `T0, 16'd540};

assign memory[247]={`LW, `T1, `T0, 16'd416};

assign memory[249]={`LW, `T1, `T0, 16'd564};

assign memory[251]={`LW, `T1, `T0, 16'd1596};

assign memory[253]={`LW, `T1, `T0, 16'd3640};

assign memory[255]={`LW, `T1, `T0, 16'd624};

assign memory[257]={`LW, `T1, `T0, 16'd3380};

assign memory[259]={`LW, `T1, `T0, 16'd2672};

assign memory[261]={`LW, `T1, `T0, 16'd820};

assign memory[263]={`LW, `T1, `T0, 16'd2496};

assign memory[265]={`LW, `T1, `T0, 16'd892};

assign memory[267]={`LW, `T1, `T0, 16'd584};

assign memory[269]={`LW, `T1, `T0, 16'd264};

assign memory[271]={`LW, `T1, `T0, 16'd156};

assign memory[273]={`LW, `T1, `T0, 16'd412};

assign memory[275]={`LW, `T1, `T0, 16'd2484};

assign memory[277]={`LW, `T1, `T0, 16'd3192};

assign memory[279]={`LW, `T1, `T0, 16'd64};

assign memory[281]={`LW, `T1, `T0, 16'd3888};

assign memory[283]={`LW, `T1, `T0, 16'd1944};

assign memory[285]={`LW, `T1, `T0, 16'd1540};

assign memory[287]={`LW, `T1, `T0, 16'd1188};

assign memory[289]={`LW, `T1, `T0, 16'd2712};

assign memory[291]={`LW, `T1, `T0, 16'd2204};

assign memory[293]={`LW, `T1, `T0, 16'd2136};

assign memory[295]={`LW, `T1, `T0, 16'd2808};

assign memory[297]={`LW, `T1, `T0, 16'd3340};

assign memory[299]={`LW, `T1, `T0, 16'd1100};

assign memory[301]={`LW, `T1, `T0, 16'd2272};

assign memory[303]={`LW, `T1, `T0, 16'd3796};

assign memory[305]={`LW, `T1, `T0, 16'd1840};

assign memory[307]={`LW, `T1, `T0, 16'd268};

assign memory[309]={`LW, `T1, `T0, 16'd76};

assign memory[311]={`LW, `T1, `T0, 16'd476};

assign memory[313]={`LW, `T1, `T0, 16'd2476};

assign memory[315]={`LW, `T1, `T0, 16'd1272};

assign memory[317]={`LW, `T1, `T0, 16'd3748};

assign memory[319]={`LW, `T1, `T0, 16'd3264};

assign memory[321]={`LW, `T1, `T0, 16'd1564};

assign memory[323]={`LW, `T1, `T0, 16'd1440};

assign memory[325]={`LW, `T1, `T0, 16'd3152};

assign memory[327]={`LW, `T1, `T0, 16'd496};

assign memory[329]={`LW, `T1, `T0, 16'd3252};

assign memory[331]={`LW, `T1, `T0, 16'd3384};

assign memory[333]={`LW, `T1, `T0, 16'd256};

assign memory[335]={`LW, `T1, `T0, 16'd3556};

assign memory[337]={`LW, `T1, `T0, 16'd1824};

assign memory[339]={`LW, `T1, `T0, 16'd1412};

assign memory[341]={`LW, `T1, `T0, 16'd3152};

assign memory[343]={`LW, `T1, `T0, 16'd948};

assign memory[345]={`LW, `T1, `T0, 16'd2204};

assign memory[347]={`LW, `T1, `T0, 16'd2708};

assign memory[349]={`LW, `T1, `T0, 16'd2512};

assign memory[351]={`LW, `T1, `T0, 16'd2316};

assign memory[353]={`LW, `T1, `T0, 16'd1156};

assign memory[355]={`LW, `T1, `T0, 16'd2604};

assign memory[357]={`LW, `T1, `T0, 16'd2504};

assign memory[359]={`LW, `T1, `T0, 16'd2072};

assign memory[361]={`LW, `T1, `T0, 16'd2412};

assign memory[363]={`LW, `T1, `T0, 16'd1648};

assign memory[365]={`LW, `T1, `T0, 16'd3704};

assign memory[367]={`LW, `T1, `T0, 16'd252};

assign memory[369]={`LW, `T1, `T0, 16'd2008};

assign memory[371]={`LW, `T1, `T0, 16'd340};

assign memory[373]={`LW, `T1, `T0, 16'd1596};

assign memory[375]={`LW, `T1, `T0, 16'd3988};

assign memory[377]={`LW, `T1, `T0, 16'd1028};

assign memory[379]={`LW, `T1, `T0, 16'd3860};

assign memory[381]={`LW, `T1, `T0, 16'd496};

assign memory[383]={`LW, `T1, `T0, 16'd2220};

assign memory[385]={`LW, `T1, `T0, 16'd3132};

assign memory[387]={`LW, `T1, `T0, 16'd3276};

assign memory[389]={`LW, `T1, `T0, 16'd3376};

assign memory[391]={`LW, `T1, `T0, 16'd768};

assign memory[393]={`LW, `T1, `T0, 16'd2084};

assign memory[395]={`LW, `T1, `T0, 16'd892};

assign memory[397]={`LW, `T1, `T0, 16'd2588};

assign memory[399]={`LW, `T1, `T0, 16'd3404};

assign memory[401]={`LW, `T1, `T0, 16'd1948};

assign memory[403]={`LW, `T1, `T0, 16'd3380};

assign memory[405]={`LW, `T1, `T0, 16'd124};

assign memory[407]={`LW, `T1, `T0, 16'd1444};

assign memory[409]={`LW, `T1, `T0, 16'd116};

assign memory[411]={`LW, `T1, `T0, 16'd1808};

assign memory[413]={`LW, `T1, `T0, 16'd560};

assign memory[415]={`LW, `T1, `T0, 16'd3472};

assign memory[417]={`LW, `T1, `T0, 16'd1720};

assign memory[419]={`LW, `T1, `T0, 16'd568};

assign memory[421]={`LW, `T1, `T0, 16'd388};

assign memory[423]={`LW, `T1, `T0, 16'd1472};

assign memory[425]={`LW, `T1, `T0, 16'd2548};

assign memory[427]={`LW, `T1, `T0, 16'd3492};

assign memory[429]={`LW, `T1, `T0, 16'd108};

assign memory[431]={`LW, `T1, `T0, 16'd800};

assign memory[433]={`LW, `T1, `T0, 16'd2328};

assign memory[435]={`LW, `T1, `T0, 16'd640};

assign memory[437]={`LW, `T1, `T0, 16'd1076};

assign memory[439]={`LW, `T1, `T0, 16'd464};

assign memory[441]={`LW, `T1, `T0, 16'd2412};

assign memory[443]={`LW, `T1, `T0, 16'd1752};

assign memory[445]={`LW, `T1, `T0, 16'd528};

assign memory[447]={`LW, `T1, `T0, 16'd2576};

assign memory[449]={`LW, `T1, `T0, 16'd2944};

assign memory[451]={`LW, `T1, `T0, 16'd3192};

assign memory[453]={`LW, `T1, `T0, 16'd3776};

assign memory[455]={`LW, `T1, `T0, 16'd3072};

assign memory[457]={`LW, `T1, `T0, 16'd4028};

assign memory[459]={`LW, `T1, `T0, 16'd2404};

assign memory[461]={`LW, `T1, `T0, 16'd3240};

assign memory[463]={`LW, `T1, `T0, 16'd244};

assign memory[465]={`LW, `T1, `T0, 16'd3784};

assign memory[467]={`LW, `T1, `T0, 16'd2016};

assign memory[469]={`LW, `T1, `T0, 16'd3512};

assign memory[471]={`LW, `T1, `T0, 16'd3052};

assign memory[473]={`LW, `T1, `T0, 16'd2160};

assign memory[475]={`LW, `T1, `T0, 16'd3568};

assign memory[477]={`LW, `T1, `T0, 16'd456};

assign memory[479]={`LW, `T1, `T0, 16'd892};

assign memory[481]={`LW, `T1, `T0, 16'd3764};

assign memory[483]={`LW, `T1, `T0, 16'd4076};

assign memory[485]={`LW, `T1, `T0, 16'd3552};

assign memory[487]={`LW, `T1, `T0, 16'd564};

assign memory[489]={`LW, `T1, `T0, 16'd3924};

assign memory[491]={`LW, `T1, `T0, 16'd1984};

assign memory[493]={`LW, `T1, `T0, 16'd2512};

assign memory[495]={`LW, `T1, `T0, 16'd2140};

assign memory[497]={`LW, `T1, `T0, 16'd160};

assign memory[499]={`LW, `T1, `T0, 16'd1384};

assign memory[501]={`LW, `T1, `T0, 16'd80};

assign memory[503]={`LW, `T1, `T0, 16'd1656};

assign memory[505]={`LW, `T1, `T0, 16'd1356};

assign memory[507]={`LW, `T1, `T0, 16'd2252};

assign memory[509]={`LW, `T1, `T0, 16'd3824};

assign memory[511]={`LW, `T1, `T0, 16'd3988};


endmodule
